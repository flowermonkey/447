////
//// Internal signal constants
////

// ALU
`define ALU_ADD      4'b0000
`define ALU_SUB      4'b0001
`define ALU_AND      4'b0010
`define ALU_OR       4'b0011
`define ALU_NOR      4'b0100
`define ALU_XOR      4'b0101
