////
//// Internal signal constants
////

// ALU
`define ALU_ADD      4'b0000
`define ALU_SUB      4'b0001
`define ALU_AND      4'b0010
`define ALU_OR       4'b0011
`define ALU_NOR      4'b0100
`define ALU_XOR      4'b0101
`define ALU_SLT      4'b0110
`define ALU_SLTU     4'b0111
`define MEM_BYTE     3'b000
`define MEM_U_BYTE   3'b100
`define MEM_HALF     3'b001
`define MEM_U_HALF   3'b101
`define MEM_WORD     3'b010
